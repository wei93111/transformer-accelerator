module matrix_mult (
    input  i_clk,
    input  i_rst_n,

);

endmodule
