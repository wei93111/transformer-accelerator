`ifndef DEFINE_VH
`define DEFINE_VH

    // operation modes
    `define INT8     0
    `define INT4     1
    `define INT4_VSQ 2
    
`endif