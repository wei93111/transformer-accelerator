`include "define.vh"

module gemm (
    input        i_clk,
    input        i_rst_n,
    input  [1:0] i_mode  

);



endmodule
