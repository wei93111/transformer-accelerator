`include "define.vh"

module mm (
    input  i_clk,
    input  i_rst_n,
    input  [1:0] i_mode,
    input 

);

endmodule
